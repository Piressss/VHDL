---------------------------------------------------------------------
-- @Author: Felipe Pires
-- @Date  : 27/12/2018
-- @Lib   : BASE LIB
-- @Code  : BASE_LIB_PKG
---------------------------------------------------------------------
package base_lib_pkg is

    -- TYPE VECTORS
    type bit1vec_t is std_logic_vector(0 downto 0);

end base_lib_pkg;
 
